* Simulación de mosfet como amplificador

*---------- DMWS120H100SM4 Spice Model ----------
.SUBCKT DMWS120H100SM4 10 20 30 
* TERMINALS : D G S
* MODEL FORMAT : SPICE3
* Editor : JAY
M1 1 2 3 3 NMOS L = 1E-06 W = 1E-06 
RD 10 1 0.055 
RS 30 3 1E-06 
RG 20 2 8.26 
CGS 2 3 1.53E-09 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1 VFB 1 
CGD 13 14 1.323E-09 
R1 13 0 1 
D1 12 13 DLIM 
DDG 15 14 DCGD 
R2 12 15 1 
D2 15 0 DLIM 
DSD 3 10 DSUB 
.MODEL NMOS NMOS LEVEL = 3 VMAX = 1E+05 ETA = 0 VTO = 4.8 TOX = 1E-07 NSUB = 8.792E+15 KP = 4.5 U0 = 100 KAPPA = 0.2 IS = 0 
.MODEL DCGD D CJO = 6E-10 VJ = 0.6 M = 0.6913 
.MODEL DSUB D IS = 3E-07 N = 8.6 RS = 0.03 BV = 1377 CJO = 1.5E-09 VJ = 0.9 M = 0.5 XTI = 0 TT = 4.94E-09 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes Spice Model v1.2 Last Revised 2023/01/10
*The model is an approximation of the device, and it may not show the true device performance under all conditions.
*The model only guarantees the accuracy of the key parameters (Ron, VSD, IDSS, Ciss, Coss, Crss, and Trr) at 25 degC in the current data sheet.

VGS Vg 0 DC 6  
X1  Vd Vg 0 DMWS120H100SM4 
*R1  Vdd VR1 2.0K
Vmean Vdd Vd DC 0
VDS Vdd 0 DC 21


*Pto. de Operación
.control
    *VOLCADO FICHERO .CIR ANALIZADO SINTACTICAMENTE
    listing > bjt.lst
    *ANALISIS PUNTO DE OPERACION
    op
    rusage everything > op.ope
    print V(Vd) V(Vg) > op.txt
    display > op.var
.endc

*Plotear Gráficas

* Obtener el valor de Vth
.control
    DC VGS 0 7 0.002
    *gnuplot graf_Ivds i(Vtest)
.endc

.control
    DC VGS 0 7 0.001
    *gnuplot graf_Ivgs -i(VGS)
.endc

* Región de Corte (𝑉𝐺𝑆<𝑉𝑡ℎ)
.control
    DC VGS 0 5 0.001 
    *gnuplot graf_R_Corte -i(VDS)
.endc


* Región de Lineal (𝑉𝐺𝑆>𝑉𝑡ℎ y VDS< VGS−Vth)

.control
    DC VDS 0 5 0.01 VGS 0 6 0.5
    gnuplot graf_R_Lineal -i(Vmean)
.endc

* Región de Saturación (VDS > VGS−Vth)

.control
    DC VDS 0 40 0.01 VGS 0 1 0.5 
    *gnuplot graf_IVds1 -i(VDS)
.endc

.end
