* SIMULATION DE-MOSFET NMOS MODEL

VGS Vg 0 DC 6  
M1  Vd Vg 0 0 IXTT20N50D 
*R1  Vdd Vd 1
VDS Vd 0 DC 21

*---------- IXTT20N50D Spice Model ----------

* IXTT20N50D Depletion NMOS model
* updated using Model Editor release 10.0.0 on 04/03/06 at 12:17
* The Model Editor is a PSpice product.
.MODEL IXTT20N50D NMOS M
+ LEVEL=3
+ L=2.0000E-6
+ W=5.5000
+ KP=1.0446E-6
+ RS=1.0000E-3
+ RD=.22202
+ VTO=-1
+ RDS=20.000E6
+ TOX=2.0000E-6
+ CGSO=6.3E-9
+ CGDO=82E-12
+ CBD=4.8729E-9
+ MJ=1.5000
+ PB=2.6055
+ RG=10.000E-3
+ IS=25E-6
+ N=2.0283
+ RB=1.0000E-9
+ GAMMA=0
+ KAPPA=0

*Pto. de Operación
.control
    *VOLCADO FICHERO .CIR ANALIZADO SINTACTICAMENTE
    listing > de-mosfet.lst
    *ANALISIS PUNTO DE OPERACION
    op
    rusage everything > op_de-mosfet.ope
    print V(Vd) V(Vg) > op_de-mosfet.txt
    display > op_de-mosfet.var
.endc

*Plotear Gráficas

****** T2.2 *****

* Región de Corte (𝑉𝐺𝑆<𝑉𝑡ℎ)
* - ID vs VGS (Verificar el valor de Vth)
.control
    DC VGS -2 0.5 0.01
    gnuplot graf_Id_vs_VGS_de-mosfet -i(VDS)
.endc

* Región de Lineal (𝑉𝐺𝑆>𝑉𝑡ℎ y VDS<VGS−Vth)
* - Id VS VDS
.control
    DC VDS 0 10 0.05 VGS -2 2 0.5
    gnuplot graf_Id_vs_VDS_de-mosfet -i(VDS)
.endc

* Región de Saturación (VDS > VGS−Vth)
.control
    DC VDS 0 40 0.1 VGS -1 2 0.5 
    gnuplot graf_Saturacion_de-mosfet -i(VDS)
.endc

.end
